// Global symbols and constants for the Pong game

`define BALL_SIZE 8 //in reaity 9 as we used <= instead of = for drawing, but didn't change the rest of the code, as not necessary
`define BALL_CENTER_OFFSET 4
`define BALL_COLOR 3'b111

`define PLAYER_HEIGHT 60
`define HALF_PLAYER_HEIGHT 30
`define PLAYER_WIDTH 12

`define FRAME_WIDTH 640
`define HALF_FRAME_WIDTH 320
`define FRAME_HEIGHT 480

`define INITIAL_BALL_X_POS 318
`define INITIAL_BALL_Y_POS 238
`define INITIAL_PLAYER_Y_POS 210

`define PLAYER_1_X_POS 13
`define PLAYER_2_X_POS 615

`define PLAYER_1_COLOR 3'b011
`define PLAYER_2_COLOR 3'b100

`define DEFAULT_PLAYER_SPEED 3

`define INITIAL_BALL_DIRECTION 0

`define COLLISION_OFFSET 4

`define CORNER_HIT_ZONE_SIZE 4
`define HIT_ZONE_1    0
`define HIT_ZONE_2   11
`define HIT_ZONE_3   23
`define HIT_ZONE_4   35
`define HIT_ZONE_5   47
`define HIT_ZONE_MAX 59

`define VERTICAL_SCORE_OFFSET 14
`define HORIZONTAL_SCORE_OFFSET 160
`define SCORE_WIDTH 16

`define WIN_TEXT_PLAYER_1_X_POS 60
`define WIN_TEXT_PLAYER_2_X_POS 520
`define WIN_TEXT_Y_POS 194

`define MENU_TEXT_X_POS 100  // z. B. Position nach Bedarf
`define MENU_TEXT_Y_POS 50
