
module rotary_encoder (
    input wire clk,
    input wire in_a,
    input wire in_b,
    input wire switch,

    output wire up,
    output wire down,
    output wire button
);
    reg a_up_first = 0;
    reg b_up_first = 0;

    reg up_r = 0;
    reg down_r = 0;
    assign up = up_r;
    assign down = down_r;

    always @(posedge clk) begin
        if (!a_up_first && !b_up_first) begin
            if (in_a) begin
                a_up_first <= 1;
            end else if (in_b) begin
                b_up_first <= 1;
            end
            up_r <= 0;
            down_r <= 0;
        end else if (a_up_first) begin
            if (in_b) begin
                up_r <= 1;
                a_up_first <= 0;
                b_up_first <= 0;
            end else begin
                up_r <= 0;
            end
        end else if (b_up_first) begin
            if (in_a) begin
                down_r <= 1;
                a_up_first <= 0;
                b_up_first <= 0;
            end else begin
                down_r <= 0;
            end
        end
    end

endmodule
