
module animation (
    input wire BALL_CLOCK,
    input wire goal_player_1,
    input wire goal_player_2,
    input wire win_player_1,
    input wire win_player_2,

    output wire[7:0] led
);
    reg goal_1_animation_triggered = 0;
    reg goal_2_animation_triggered = 0;
    reg win_1_animation_triggered = 0;
    reg win_2_animation_triggered = 0;

    reg[7:0] led_r;
    assign led = led_r;

    reg[1:0] repetitions = 0;

    reg[1:0] delay = 2'b11;

    always @(posedge BALL_CLOCK) begin
        if (goal_1_animation_triggered && (repetitions != 2'b0)) begin
            casez ({delay, led_r})
                10'b11_????????: delay <= delay - 1;
                10'b10_????????: delay <= delay - 1;
                10'b01_????????: delay <= delay - 1;

                10'b00_00000000: led_r <= 8'b10000000;
                10'b00_10000000: led_r <= 8'b01000000;
                10'b00_01000000: led_r <= 8'b00100000;
                10'b00_00100000: led_r <= 8'b00010000;
                10'b00_00010000: led_r <= 8'b00001000;
                10'b00_00001000: led_r <= 8'b00000100;
                10'b00_00000100: led_r <= 8'b00000010;
                10'b00_00000010: led_r <= 8'b00000001;
                10'b00_00000001: begin
                    led_r <= 8'b00000000;
                    repetitions <= repetitions - 1;
                end
                default: led_r <= 0;
            endcase

        end else if (goal_2_animation_triggered && (repetitions != 2'b0)) begin
            casez ({delay, led_r})
                10'b11_????????: delay <= delay - 1;
                10'b10_????????: delay <= delay - 1;
                10'b01_????????: delay <= delay - 1;

                10'b00_00000000: led_r <= 8'b00000001;
                10'b00_00000001: led_r <= 8'b00000010;
                10'b00_00000010: led_r <= 8'b00000100;
                10'b00_00000100: led_r <= 8'b00001000;
                10'b00_00001000: led_r <= 8'b00010000;
                10'b00_00010000: led_r <= 8'b00100000;
                10'b00_00100000: led_r <= 8'b01000000;
                10'b00_01000000: led_r <= 8'b10000000;
                10'b00_10000000: begin
                    led_r <= 8'b00000000;
                    repetitions <= repetitions - 1;
                end 
                default: led_r <= 0;
            endcase

        end else if (win_1_animation_triggered && (repetitions != 2'b0)) begin
            casez ({delay, led_r})
                10'b11_????????: delay <= delay - 1;
                10'b10_????????: delay <= delay - 1;
                10'b01_????????: delay <= delay - 1;

                10'b00_00000000: led_r <= 8'b10000001;
                10'b00_10000001: led_r <= 8'b01000010;
                10'b00_01000010: led_r <= 8'b00100100;
                10'b00_00100100: led_r <= 8'b00011000;
                10'b00_00011000: led_r <= 8'b00111000;
                10'b00_00111000: led_r <= 8'b01111000;
                10'b00_01111000: led_r <= 8'b11111000;
                10'b00_11111000: begin
                    led_r <= 8'b00000000;
                    repetitions <= repetitions - 1;
                end
                default: led_r <= 0;
            endcase

        end else if (win_2_animation_triggered && (repetitions != 2'b0)) begin
            casez ({delay, led_r})
                10'b11_????????: delay <= delay - 1;
                10'b10_????????: delay <= delay - 1;
                10'b01_????????: delay <= delay - 1;

                10'b00_00000000: led_r <= 8'b10000001;
                10'b00_10000001: led_r <= 8'b01000010;
                10'b00_01000010: led_r <= 8'b00100100;
                10'b00_00100100: led_r <= 8'b00011000;
                10'b00_00011000: led_r <= 8'b00011100;
                10'b00_00011100: led_r <= 8'b00011110;
                10'b00_00011110: led_r <= 8'b00011111;
                10'b00_00011111: begin
                    led_r <= 8'b00000000;
                    repetitions <= repetitions - 1;
                end
                default: led_r <= 0;
            endcase

        end else begin
            led_r <= 8'b0;
            if (win_player_1) begin
                win_1_animation_triggered <= 1;
                win_2_animation_triggered <= 0;
                goal_1_animation_triggered <= 0;
                goal_2_animation_triggered <= 0;

            end if (win_player_2) begin
                win_1_animation_triggered <= 0;
                win_2_animation_triggered <= 1;
                goal_1_animation_triggered <= 0;
                goal_2_animation_triggered <= 0;

            end if (goal_player_1) begin
                win_1_animation_triggered <= 0;
                win_2_animation_triggered <= 0;
                goal_1_animation_triggered <= 1;
                goal_2_animation_triggered <= 0;

            end if (goal_player_2) begin
                win_1_animation_triggered <= 0;
                win_2_animation_triggered <= 0;
                goal_1_animation_triggered <= 0;
                goal_2_animation_triggered <= 1;
            end

            if (win_player_1 || win_player_2 || goal_player_1 || goal_player_2) begin
                repetitions <= 2'b11;
            end
        end
    end

endmodule
